this is not an entity 
